`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   22:08:52 03/29/2021
// Design Name:   ppl
// Module Name:   D:/Code/WebISE/lab92Ryan/ppl/bench.v
// Project Name:  ppl
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: ppl
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module bench;

	// Inputs
	reg clk;	
	reg downloading;
	reg [1:0] flag;
	reg [31:0] instrc;
	reg rst;
	reg detect;
	reg [9:0] det_addr;
	wire [31:0] det_data;

	// Instantiate the Unit Under Test (UUT)
	cmt uut (
		.clk(clk), 		
		.downloading(downloading),
		.flag(flag),
		.instrc(instrc),
		.rst(rst),
		.detect(detect),
		.det_addr(det_addr),
		.det_data(det_data)
	);

	initial begin
		// Initialize Inputs
		clk = 1'b0;		
		downloading = 1'b0;
		instrc = 32'h00000000;
		flag=2'b00;
		rst=1'b0;
		detect=1'b0;
		det_addr=10'b0000000000;
		#25
		// Wait 100 ns for global reset to finish
//////////////////////////////////////////////thread0///////////////////////////////////////
		instrc=32'hfd010113;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h02812623;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h03010413;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00100793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfcf42823;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00200793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfcf42a23;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00300793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfcf42c23;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00400793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfcf42e23;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00500793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfef42023;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe042623;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h0c80006f;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe042423;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h0a00006f;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040713;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f707b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe07a703;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00178793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040693;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f687b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe07a783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h06f75263;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040713;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f707b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe07a783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfef42223;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00178793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040713;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f707b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe07a703;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040693;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f687b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfee7a023;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00178793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040713;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f707b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe442703;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfee7a023;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00178793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfef42423;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00400713;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfec42783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h40f707b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842703;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hf4f74ae3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfec42783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00178793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfef42623;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfec42703;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00300793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hf2e7dae3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00000013;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00000013;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h02c12403;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h03010113;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00008067;
		downloading=1'b0;
		#50
		downloading=1'b1;		
		#50			
	//////////////////////////////////////thread1///////////////////////////////////////////
		flag=2'b01;
		instrc=32'hfd010113;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h02812623;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h03010413;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00100793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfcf42823;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00200793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfcf42a23;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00300793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfcf42c23;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00400793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfcf42e23;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00500793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfef42023;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe042623;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h0c80006f;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe042423;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h0a00006f;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040713;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f707b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe07a703;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00178793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040693;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f687b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe07a783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h06f75263;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040713;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f707b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe07a783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfef42223;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00178793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040713;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f707b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe07a703;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040693;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f687b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfee7a023;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00178793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040713;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f707b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe442703;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfee7a023;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00178793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfef42423;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00400713;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfec42783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h40f707b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842703;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hf4f74ae3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfec42783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00178793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfef42623;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfec42703;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00300793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hf2e7dae3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00000013;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00000013;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h02c12403;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h03010113;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00008067;
		downloading=1'b0;
		#50
		downloading=1'b1;		
		#50			
	//////////////////////////////////////thread2///////////////////////////////////////////
		flag=2'b10;
		instrc=32'hfd010113;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h02812623;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h03010413;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00100793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfcf42823;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00200793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfcf42a23;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00300793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfcf42c23;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00400793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfcf42e23;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00500793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfef42023;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe042623;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h0c80006f;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe042423;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h0a00006f;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040713;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f707b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe07a703;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00178793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040693;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f687b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe07a783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h06f75263;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040713;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f707b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe07a783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfef42223;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00178793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040713;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f707b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe07a703;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040693;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f687b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfee7a023;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00178793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040713;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f707b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe442703;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfee7a023;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00178793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfef42423;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00400713;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfec42783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h40f707b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842703;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hf4f74ae3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfec42783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00178793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfef42623;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfec42703;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00300793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hf2e7dae3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00000013;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00000013;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h02c12403;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h03010113;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00008067;
		downloading=1'b0;
		#50
		downloading=1'b1;		
		#50	
		///////////////////////////////////////thread3///////////////////////////////////////////
		flag=2'b11;
		instrc=32'hfd010113;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h02812623;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h03010413;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00100793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfcf42823;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00200793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfcf42a23;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00300793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfcf42c23;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00400793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfcf42e23;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00500793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfef42023;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe042623;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h0c80006f;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe042423;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h0a00006f;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040713;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f707b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe07a703;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00178793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040693;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f687b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe07a783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h06f75263;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040713;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f707b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe07a783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfef42223;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00178793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040713;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f707b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe07a703;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040693;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f687b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfee7a023;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00178793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00279793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hff040713;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00f707b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe442703;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfee7a023;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00178793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfef42423;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00400713;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfec42783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h40f707b3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfe842703;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hf4f74ae3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfec42783;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00178793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfef42623;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hfec42703;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00300793;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'hf2e7dae3;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00000013;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00000013;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h02c12403;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h03010113;
		downloading=1'b0;
		#50
		downloading=1'b1;
		#50
		instrc=32'h00008067;
		downloading=1'b0;
		#50
		downloading=1'b1;		
		#50	
		downloading=1'b0;
		#25
		rst=1'b1;
		#900000
		detect=1'b1;
		det_addr=10'b1111110100;
		#50
		$stop;
		
		
		// Add stimulus here

	end
	
	always
	begin
		#25
			clk=~clk;
   end
	
	
endmodule

